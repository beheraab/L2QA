************************************************************************
* auCdl Netlist:
* 
* Library Name:  flat_schematic_lib
* Top Cell Name: i0minv000aa1n02x5
* View Name:     schematic
* Netlisted on:  Jul 18 22:35:06 2021
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA



*.EXPAND_ON_M_FACTOR

************************************************************************
* Library Name: flat_schematic_lib
* Cell Name:    i0minv000aa1n02x5
* View Name:    schematic
************************************************************************

.SUBCKT i0minv000aa1n02x5 a o1 vcc vssx
*.PININFO a:I o1:O vcc:B vssx:B
Mg101.qna.mn2 o1 a vssx vssx nhpaulvt W=2.0 L=14n m=1 lvsExactMatch=1
Mg101.qpa.mp2 o1 a vcc vcc phpaulvt W=2.0 L=14n m=1 lvsExactMatch=1
.ENDS
